entity mux is
    port (
        I : in std_logic_vector (3 downto 0); 
        SEL : in std_logic_vector (1 downto 0); 
        Y : out std_logic 
    );
end entity mux;

architecture behav_mux of mux is 
begin 

    

end architecture behav_mux; 